// comment
/* anot
ther
com
ment*/

/*yikes*/c/*a*/las/**/s test; // jfjfj
endclas/*jabs*/s
