`include "task0.svh"
`include "task1.svh"
`include "task2.svh"
`include "task3.svh"
`include "task4.svh"
`include "task5.svh"
`include "task6.svh"
`include "task7.svh"
