`define WIDTH 1
