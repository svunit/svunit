automatic function int unsigned factorial(int unsigned n);
  return 0;
endfunction
