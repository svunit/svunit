interface static test_if2();
endinterface
