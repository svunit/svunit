test-xyz.abc-
