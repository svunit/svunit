module dut;
  module_in_my_filelist m();
endmodule
