`include "write.svh"
