class queue;
endclass
