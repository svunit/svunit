/**
 * Extracts the full name of a test from the return value of $typename.
 *
 * The return value of $typename varies wildly across simulators.
 */
class full_name_extraction;

  function string get_full_name(string dollar_typename);
    // TODO Implement
  endfunction

endclass
