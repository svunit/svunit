class testcase extends svunit_testcase;

  function new(string name);
    super.new(name);
  endfunction

endclass
