package factorial;

  function automatic int unsigned factorial(int unsigned n);
    return 1;
  endfunction

endpackage
