library verilog;
use verilog.vl_types.all;
entity \__home_njohnson_work_svunit_code_test_svunit_base_0b_testsuite_sv_unit\ is
end \__home_njohnson_work_svunit_code_test_svunit_base_0b_testsuite_sv_unit\;
