interface dut;
endinterface
