module automatic test_automatic();
endmodule
