`ifndef SVUNIT_TYPES
`define SVUNIT_TYPES

  /*
    Enum: results_t
    enumerated type containing PASS/FAIL
  */
  typedef enum {PASS=1, FAIL=0}  results_t;


  /*
    Enum: boolean_t
    enumerated type containing TRUE/FALSE
  */
  typedef enum {TRUE=1, FALSE=0} boolean_t;

`endif
