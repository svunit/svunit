class test2;
endclass
