class dut;
endclass
