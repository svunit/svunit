class subdir1a;
endclass
