package a_pkg;
  class a_class;
  endclass
endpackage
