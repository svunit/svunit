module dut;
  wire a, b, c;
  vhd_e vhd_e(a, b, c);
endmodule
