module another_filelist_module();
  yet_another_module yam();
endmodule
