class stack;
endclass
