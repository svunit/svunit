class queue;

  function int unsigned size();
    return 0;
  endfunction


  function void push(int unsigned elem);
  endfunction

endclass
