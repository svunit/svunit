class test0;
endclass

class test1;
endclass
