package data_structures;

  `include "queue.svh"
  `include "stack.svh"

endpackage
