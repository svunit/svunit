class subdir1;
endclass
