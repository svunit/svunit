module module_in_my_filelist;
  another_filelist_module a();
endmodule
