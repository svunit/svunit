module svunit_main;

  // initial
  //   svunit::run_all_tests();

endmodule
