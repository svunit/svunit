library verilog;
use verilog.vl_types.all;
entity dut_unit_test is
end dut_unit_test;
