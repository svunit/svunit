package test_data_structures;

  import data_structures::*;

  `include "test_queue.svh"
  `include "test_stack.svh"

endpackage
