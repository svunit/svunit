class test_queue;

  // TODO Add tests for `queue`

endclass
