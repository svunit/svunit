class test0;
endclass

class test1;
endclass

virtual class test2;
endclass
