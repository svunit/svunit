module dut;
endmodule
