// The current testcase that is being executed.
svunit_testcase current_tc;
