class test_stack;

  // TODO Add tests for `stack`

endclass
