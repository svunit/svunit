class test0;
endclass
