module my_and_module
(
  input a,
  input b,
  output wire ab
);

assign ab = a && b;

endmodule
