//###########################################################################
//
//  Copyright 2024 The SVUnit Authors.
//
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
//
//###########################################################################

/*
  Base class for tests defined using the `SVTEST macro
*/
virtual class svunit_test extends svunit_base;

  function new(string name);
    super.new(name);
  endfunction


  pure virtual task unit_test_setup();
  pure virtual task run();
  pure virtual task unit_test_teardown();

endclass
