// comment
/* anot
ther
com
ment*/

/*//
//*/
/*//*/
/*yikes*/c/*a*/las/**/s virtual_test; // jfjfj
endclas/*jabs*/s
