/**
 * A dummy type that can be used in places where a type is required by the compiler, but the type
 * is irrelevant. One such place is as a default for type parameters, because some simulators
 * do not allow parameters without default values.
 */
class dummy;

  // Intentionally empty

endclass
