package factorial;

  function automatic int unsigned factorial(int unsigned n);
    return 0;
  endfunction

endpackage
