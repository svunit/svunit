module another_filelist_module();
endmodule
