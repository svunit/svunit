class stack;

  function int unsigned size();
    return 0;
  endfunction

endclass
