class subdir0;
endclass
