library verilog;
use verilog.vl_types.all;
entity svunit_pkg is
end svunit_pkg;
