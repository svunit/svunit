`ifndef __AMBA_XACTION__
`define __AMBA_XACTION__

class amba_xaction extends vmm_data;
endclass


`endif
