module static test_static();
endmodule
