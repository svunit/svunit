//###########################################################################
//
//  Copyright 2011 The SVUnit Authors.
//
//  Licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing, software
//  distributed under the License is distributed on an "AS IS" BASIS,
//  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//  See the License for the specific language governing permissions and
//  limitations under the License.
//
//###########################################################################

`ifndef SVUNIT_TYPES
`define SVUNIT_TYPES

  /*
    Enum: results_t
    enumerated type containing PASS/FAIL
  */
  typedef enum {PASS=1, FAIL=0}  results_t;


  /*
    Enum: boolean_t
    enumerated type containing TRUE/FALSE
  */
  typedef enum {TRUE=1, FALSE=0} boolean_t;

`endif
