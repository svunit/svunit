module test();
endmodule
