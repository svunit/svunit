class test3;
endclass
