package queue;

  class queue #(type T = int);

    function void enqueue(T e);
    endfunction

  endclass

endpackage
