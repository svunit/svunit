class test_registry;

  function void register(test::builder test_builder, string full_name);
    // TODO Implement
  endfunction

endclass
