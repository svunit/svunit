interface test_if();
endinterface
