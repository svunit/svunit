package test_data_structures;

  import data_structures::*;

  `include "svunit.svh"
  `include "svunit_defines.svh"

  `include "test_queue.svh"
  `include "test_stack.svh"

endpackage
