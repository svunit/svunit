interface automatic test_if();
endinterface
