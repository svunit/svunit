test.xyz-
