module yet_another_module;
endmodule
